/*
<????? ??>
1. ?? ??
2. ?? ??
3. ??
4. ?? ??/?? ??
5. ???

wire, reg

alway @ ??
begin end? ????.
?? ??? ?? ??

test banch
timesacle ??? ????.


timescale 1ns/100ps
module Tb_AND
...



*/

module not_gate (
	input a,
	output y
);
	//wire a;		//??, ?? ??? ? ??.
	assign y=~a;

endmodule