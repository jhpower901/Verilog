`timescale 1ns/100ps
module cycle (clk, init_val_chk, x, cycle_chk);
	input wire clk;
	input wire init_val_chk;
	input wire [7:0] x;
	output reg cycle_chk;
	reg [7:0] state_1;
	reg [7:0] state_2;

	always @(init_val_chk) begin
		flag = 0;
		state_1 = 8'b0000_0000;
		state_2 = 8'b0000_0000;
	end

	always @(posedge clk) begin
		if (state_2 == x)
			flag = 1;
		else
			flag = 0;
		state_2 = state_1;
		state_1 = x;
	end
endmodule